`include "CONFIG_MACROS.v"

module UART_RX (input wire CLK,
                input wire RST,
                input wire RX_IN,
                input wire PAR_EN,
                input wire PAR_TYP,
                input wire [4:0] Prescale,

                output wire Data_Valid,
                output wire [`WIDTH-1:0] P_DATA);

    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////////// Internal Signals ///////////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////
    
    wire par_err_int;
    wire strt_glitch_int;
    wire stp_err_int;
    wire [`BIT_COUNTER_WIDTH-1:0] bit_cnt_int;
    wire [4:0] edge_cnt_int;
    wire par_chk_en_int;
    wire strt_chk_en_int;
    wire stp_chk_en_int;
    wire deser_en_int;
    wire edge_count_en_int;
    wire data_sample_en_int;
    wire sampled_bit_int;
    wire StartTransition_int;


    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////////// FSM Instantiation //////////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

    FSM FSM_Module (
    .CLK(CLK),
    .RST(RST),
    .RX_IN(RX_IN),
    .PAR_EN(PAR_EN),
    .par_err(par_err_int),
    .strt_glitch(strt_glitch_int),
    .stp_err(stp_err_int),
    .bit_cnt(bit_cnt_int),
    .edge_cnt(edge_cnt_int),
    .Prescale(Prescale),
    .StartTransition(StartTransition_int),
    .par_chk_en(par_chk_en_int),
    .strt_chk_en(strt_chk_en_int),
    .stp_chk_en(stp_chk_en_int),
    .Data_Valid(Data_Valid),
    .deser_en(deser_en_int),
    .edge_count_en(edge_count_en_int),
    .data_sample_en(data_sample_en_int)
    );

    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////// deserializer Instantiation /////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

    deserializer deser_Module (
    .deser_en(deser_en_int),
    .sampled_bit(sampled_bit_int),
    .CLK(CLK),
    .RST(RST),
    .P_DATA(P_DATA)
    );

    /////////////////////////////////////////////////////////////////////////////////////////////
    ///////////////////////////////// strt_check Instantiation //////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////
    
    strt_check strt_check_Module (
    .strt_chk_en(strt_chk_en_int),
    .sampled_bit(sampled_bit_int),
    .strt_glitch(strt_glitch_int)
    );

    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////// parity_check Instantiation /////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

    parity_check parity_check_Module (
    .CLK(CLK),
    .RST(RST),
    .par_chk_en(par_chk_en_int),
    .PAR_TYP(PAR_TYP),
    .sampled_bit(sampled_bit_int),
    .PAR_EN(PAR_EN),
    .P_DATA(P_DATA),
    .par_err(par_err_int)
    );
    
    /////////////////////////////////////////////////////////////////////////////////////////////
    ////////////////////////////////// stp_check Instantiation //////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

    stp_check stp_check_Module (
    .CLK(CLK),
    .RST(RST),
    .stp_chk_en(stp_chk_en_int),
    .sampled_bit(sampled_bit_int),
    
    .stp_err(stp_err_int)
    );

    /////////////////////////////////////////////////////////////////////////////////////////////
    ////////////////////////////// edge_bit_counter Instantiation ///////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

    edge_bit_counter edge_bit_counter_Module (
    .CLK(CLK),
    .RST(RST),
    .edge_count_en(edge_count_en_int),
    .Prescale(Prescale),
    .StartTransition(StartTransition_int),
    
    .bit_cnt(bit_cnt_int),
    .edge_cnt(edge_cnt_int)
    );

    /////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////// data_sampler Instantiation /////////////////////////////////
    /////////////////////////////////////////////////////////////////////////////////////////////

    data_sampler data_sampler_Module (
    .CLK(CLK),
    .RST(RST),
    .data_sample_en(data_sample_en_int),
    .RX_IN(RX_IN),
    
    .sampled_bit(sampled_bit_int)
    );
    
    
endmodule
